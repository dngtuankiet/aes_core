module tb_AES_GCM();

endmodule
