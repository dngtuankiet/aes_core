module AES_GCM();
endmodule
