module tb_AES_Block();
reg CLK;
reg RST;
reg EN;
reg [0:127] PTEXT;
reg VALID_PTEXT;
reg [0:255] KEY;
reg VALID_KEY;
wire [0:127] CTEXT;
wire VALID_CTEXT;
//-----------------------------------//

AES_Block AES_BLOCK(
.iClk(CLK),
.iRst_n(RST),
.iEn(EN),
.iPtext(PTEXT),
.iValid_Ptext(VALID_PTEXT),
.iKey(KEY),
.iValid_Key(VALID_KEY),
.oCtext(CTEXT),
.oValid_Ctext(VALID_CTEXT)
);

initial begin
CLK = 0;
RST = 0;
EN = 0;
PTEXT = 0;
VALID_PTEXT = 0;
KEY = 0;
VALID_KEY = 0;
end

always #5 CLK = ~CLK;

//PTEXT (ASCII): 123456789abcdefg
//CORESSPOND PTEXT: 0x31323334353637383961626364656667
//TEXT KEY (ASCII): 123456789abcdefg123456789abcdefg 
//CORESSPOND KEY: 0x3132333435363738396162636465666731323334353637383961626364656667
//CTEXT: 0xB5A10E6B334037DE03F8D25BFE7ADAAA

//PTEXT: 0x00112233445566778899aabbccddeeff
//KEY:	 0x000102030405060708090a0b0c0d0e0f101112131415161718191a1b1c1d1e1f
//CTEXT: 0x8ea2b7ca516745bfeafc49904b496089
initial begin
#30
@(posedge CLK)
RST = 1;
EN = 1;
#30
//first text
@(posedge CLK)
PTEXT = 128'h31323334353637383961626364656667;
VALID_PTEXT = 1;
KEY = 256'h3132333435363738396162636465666731323334353637383961626364656667;
VALID_KEY = 1;
@(posedge CLK)
PTEXT = 0;
VALID_PTEXT = 0;
KEY = 0;
VALID_KEY = 0;

@(posedge CLK);
@(posedge CLK);
@(posedge CLK);

//second text
@(posedge CLK)
PTEXT = 128'h00112233445566778899aabbccddeeff;
VALID_PTEXT = 1;
KEY = 256'h000102030405060708090a0b0c0d0e0f101112131415161718191a1b1c1d1e1f;
VALID_KEY = 1;
@(posedge CLK)
PTEXT = 0;
VALID_PTEXT = 0;
KEY = 0;
VALID_KEY = 0;


#30
@(posedge CLK)
#300
$finish;
end

endmodule
